library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

package sin256rom_pkg is
	type rom is array (0 to 255) of signed(15 downto 0);
	constant sin256rom : rom;
end sin256rom_pkg;

package body sin256rom_pkg is
	constant sin256rom : rom := (
		to_signed(0, 16),
		to_signed(804, 16),
		to_signed(1608, 16),
		to_signed(2410, 16),
		to_signed(3212, 16),
		to_signed(4011, 16),
		to_signed(4808, 16),
		to_signed(5602, 16),
		to_signed(6393, 16),
		to_signed(7179, 16),
		to_signed(7962, 16),
		to_signed(8739, 16),
		to_signed(9512, 16),
		to_signed(10278, 16),
		to_signed(11039, 16),
		to_signed(11793, 16),
		to_signed(12539, 16),
		to_signed(13279, 16),
		to_signed(14010, 16),
		to_signed(14732, 16),
		to_signed(15446, 16),
		to_signed(16151, 16),
		to_signed(16846, 16),
		to_signed(17530, 16),
		to_signed(18204, 16),
		to_signed(18868, 16),
		to_signed(19519, 16),
		to_signed(20159, 16),
		to_signed(20787, 16),
		to_signed(21403, 16),
		to_signed(22005, 16),
		to_signed(22594, 16),
		to_signed(23170, 16),
		to_signed(23731, 16),
		to_signed(24279, 16),
		to_signed(24811, 16),
		to_signed(25329, 16),
		to_signed(25832, 16),
		to_signed(26319, 16),
		to_signed(26790, 16),
		to_signed(27245, 16),
		to_signed(27683, 16),
		to_signed(28105, 16),
		to_signed(28510, 16),
		to_signed(28898, 16),
		to_signed(29268, 16),
		to_signed(29621, 16),
		to_signed(29956, 16),
		to_signed(30273, 16),
		to_signed(30571, 16),
		to_signed(30852, 16),
		to_signed(31113, 16),
		to_signed(31356, 16),
		to_signed(31580, 16),
		to_signed(31785, 16),
		to_signed(31971, 16),
		to_signed(32137, 16),
		to_signed(32285, 16),
		to_signed(32412, 16),
		to_signed(32521, 16),
		to_signed(32609, 16),
		to_signed(32678, 16),
		to_signed(32728, 16),
		to_signed(32757, 16),
		to_signed(32767, 16),
		to_signed(32757, 16),
		to_signed(32728, 16),
		to_signed(32678, 16),
		to_signed(32609, 16),
		to_signed(32521, 16),
		to_signed(32412, 16),
		to_signed(32285, 16),
		to_signed(32137, 16),
		to_signed(31971, 16),
		to_signed(31785, 16),
		to_signed(31580, 16),
		to_signed(31356, 16),
		to_signed(31113, 16),
		to_signed(30852, 16),
		to_signed(30571, 16),
		to_signed(30273, 16),
		to_signed(29956, 16),
		to_signed(29621, 16),
		to_signed(29268, 16),
		to_signed(28898, 16),
		to_signed(28510, 16),
		to_signed(28105, 16),
		to_signed(27683, 16),
		to_signed(27245, 16),
		to_signed(26790, 16),
		to_signed(26319, 16),
		to_signed(25832, 16),
		to_signed(25329, 16),
		to_signed(24811, 16),
		to_signed(24279, 16),
		to_signed(23731, 16),
		to_signed(23170, 16),
		to_signed(22594, 16),
		to_signed(22005, 16),
		to_signed(21403, 16),
		to_signed(20787, 16),
		to_signed(20159, 16),
		to_signed(19519, 16),
		to_signed(18868, 16),
		to_signed(18204, 16),
		to_signed(17530, 16),
		to_signed(16846, 16),
		to_signed(16151, 16),
		to_signed(15446, 16),
		to_signed(14732, 16),
		to_signed(14010, 16),
		to_signed(13279, 16),
		to_signed(12539, 16),
		to_signed(11793, 16),
		to_signed(11039, 16),
		to_signed(10278, 16),
		to_signed(9512, 16),
		to_signed(8739, 16),
		to_signed(7962, 16),
		to_signed(7179, 16),
		to_signed(6393, 16),
		to_signed(5602, 16),
		to_signed(4808, 16),
		to_signed(4011, 16),
		to_signed(3212, 16),
		to_signed(2410, 16),
		to_signed(1608, 16),
		to_signed(804, 16),
		to_signed(0, 16),
		to_signed(-804, 16),
		to_signed(-1608, 16),
		to_signed(-2410, 16),
		to_signed(-3212, 16),
		to_signed(-4011, 16),
		to_signed(-4808, 16),
		to_signed(-5602, 16),
		to_signed(-6393, 16),
		to_signed(-7179, 16),
		to_signed(-7962, 16),
		to_signed(-8739, 16),
		to_signed(-9512, 16),
		to_signed(-10278, 16),
		to_signed(-11039, 16),
		to_signed(-11793, 16),
		to_signed(-12539, 16),
		to_signed(-13279, 16),
		to_signed(-14010, 16),
		to_signed(-14732, 16),
		to_signed(-15446, 16),
		to_signed(-16151, 16),
		to_signed(-16846, 16),
		to_signed(-17530, 16),
		to_signed(-18204, 16),
		to_signed(-18868, 16),
		to_signed(-19519, 16),
		to_signed(-20159, 16),
		to_signed(-20787, 16),
		to_signed(-21403, 16),
		to_signed(-22005, 16),
		to_signed(-22594, 16),
		to_signed(-23170, 16),
		to_signed(-23731, 16),
		to_signed(-24279, 16),
		to_signed(-24811, 16),
		to_signed(-25329, 16),
		to_signed(-25832, 16),
		to_signed(-26319, 16),
		to_signed(-26790, 16),
		to_signed(-27245, 16),
		to_signed(-27683, 16),
		to_signed(-28105, 16),
		to_signed(-28510, 16),
		to_signed(-28898, 16),
		to_signed(-29268, 16),
		to_signed(-29621, 16),
		to_signed(-29956, 16),
		to_signed(-30273, 16),
		to_signed(-30571, 16),
		to_signed(-30852, 16),
		to_signed(-31113, 16),
		to_signed(-31356, 16),
		to_signed(-31580, 16),
		to_signed(-31785, 16),
		to_signed(-31971, 16),
		to_signed(-32137, 16),
		to_signed(-32285, 16),
		to_signed(-32412, 16),
		to_signed(-32521, 16),
		to_signed(-32609, 16),
		to_signed(-32678, 16),
		to_signed(-32728, 16),
		to_signed(-32757, 16),
		to_signed(-32767, 16),
		to_signed(-32757, 16),
		to_signed(-32728, 16),
		to_signed(-32678, 16),
		to_signed(-32609, 16),
		to_signed(-32521, 16),
		to_signed(-32412, 16),
		to_signed(-32285, 16),
		to_signed(-32137, 16),
		to_signed(-31971, 16),
		to_signed(-31785, 16),
		to_signed(-31580, 16),
		to_signed(-31356, 16),
		to_signed(-31113, 16),
		to_signed(-30852, 16),
		to_signed(-30571, 16),
		to_signed(-30273, 16),
		to_signed(-29956, 16),
		to_signed(-29621, 16),
		to_signed(-29268, 16),
		to_signed(-28898, 16),
		to_signed(-28510, 16),
		to_signed(-28105, 16),
		to_signed(-27683, 16),
		to_signed(-27245, 16),
		to_signed(-26790, 16),
		to_signed(-26319, 16),
		to_signed(-25832, 16),
		to_signed(-25329, 16),
		to_signed(-24811, 16),
		to_signed(-24279, 16),
		to_signed(-23731, 16),
		to_signed(-23170, 16),
		to_signed(-22594, 16),
		to_signed(-22005, 16),
		to_signed(-21403, 16),
		to_signed(-20787, 16),
		to_signed(-20159, 16),
		to_signed(-19519, 16),
		to_signed(-18868, 16),
		to_signed(-18204, 16),
		to_signed(-17530, 16),
		to_signed(-16846, 16),
		to_signed(-16151, 16),
		to_signed(-15446, 16),
		to_signed(-14732, 16),
		to_signed(-14010, 16),
		to_signed(-13279, 16),
		to_signed(-12539, 16),
		to_signed(-11793, 16),
		to_signed(-11039, 16),
		to_signed(-10278, 16),
		to_signed(-9512, 16),
		to_signed(-8739, 16),
		to_signed(-7962, 16),
		to_signed(-7179, 16),
		to_signed(-6393, 16),
		to_signed(-5602, 16),
		to_signed(-4808, 16),
		to_signed(-4011, 16),
		to_signed(-3212, 16),
		to_signed(-2410, 16),
		to_signed(-1608, 16),
		to_signed(-804, 16));
end package body sin256rom_pkg;
